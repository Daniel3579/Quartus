library verilog;
use verilog.vl_types.all;
entity labthirdthird_vlg_vec_tst is
end labthirdthird_vlg_vec_tst;
