library verilog;
use verilog.vl_types.all;
entity labthirdthird is
    port(
        a               : in     vl_logic;
        a1              : in     vl_logic;
        b               : in     vl_logic;
        b1              : in     vl_logic;
        k               : in     vl_logic;
        z               : in     vl_logic;
        p0              : out    vl_logic;
        p               : out    vl_logic;
        s1              : out    vl_logic;
        s               : out    vl_logic
    );
end labthirdthird;
