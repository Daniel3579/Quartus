library verilog;
use verilog.vl_types.all;
entity labthirdsecond_vlg_vec_tst is
end labthirdsecond_vlg_vec_tst;
