library verilog;
use verilog.vl_types.all;
entity labthirdsecond is
    port(
        S1              : out    vl_logic;
        A               : in     vl_logic;
        B               : in     vl_logic;
        Z               : in     vl_logic;
        S2              : out    vl_logic;
        A1              : in     vl_logic;
        B1              : in     vl_logic;
        K               : in     vl_logic;
        P               : out    vl_logic
    );
end labthirdsecond;
