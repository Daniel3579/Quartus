library verilog;
use verilog.vl_types.all;
entity labfirstsecond_vlg_vec_tst is
end labfirstsecond_vlg_vec_tst;
