library verilog;
use verilog.vl_types.all;
entity labthirdthird_vlg_sample_tst is
    port(
        a               : in     vl_logic;
        a1              : in     vl_logic;
        b               : in     vl_logic;
        b1              : in     vl_logic;
        k               : in     vl_logic;
        z               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end labthirdthird_vlg_sample_tst;
