library verilog;
use verilog.vl_types.all;
entity labfourth_vlg_vec_tst is
end labfourth_vlg_vec_tst;
