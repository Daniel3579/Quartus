library verilog;
use verilog.vl_types.all;
entity labthirdfirst_vlg_vec_tst is
end labthirdfirst_vlg_vec_tst;
