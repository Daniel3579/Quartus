library verilog;
use verilog.vl_types.all;
entity labthirdthird_vlg_check_tst is
    port(
        p               : in     vl_logic;
        p0              : in     vl_logic;
        s               : in     vl_logic;
        s1              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end labthirdthird_vlg_check_tst;
