library verilog;
use verilog.vl_types.all;
entity labthirdfirst_vlg_check_tst is
    port(
        P               : in     vl_logic;
        S               : in     vl_logic;
        S1              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end labthirdfirst_vlg_check_tst;
