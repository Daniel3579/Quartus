library verilog;
use verilog.vl_types.all;
entity labfourthsecond_vlg_vec_tst is
end labfourthsecond_vlg_vec_tst;
