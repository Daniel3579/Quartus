library verilog;
use verilog.vl_types.all;
entity labfirstfirst_vlg_vec_tst is
end labfirstfirst_vlg_vec_tst;
